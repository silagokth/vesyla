`define dummy_impl _fsahpf8ao5p
`define dummy_impl_pkg _fsahpf8ao5p_pkg


package _fsahpf8ao5p_pkg;
    parameter RESOURCE_INSTR_WIDTH = 27;
endpackage

module _fsahpf8ao5p
import _fsahpf8ao5p_pkg::*;
(
    input  logic clk_0,
    input  logic rst_n_0,
    input  logic instr_en_0,
    input  logic [RESOURCE_INSTR_WIDTH-1:0] instr_0,
    input  logic activate_0
);
endmodule
