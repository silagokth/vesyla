`define dummy_impl2 _fsahpf8ao5p
`define dummy_impl2_pkg _fsahpf8ao5p_pkg

